library verilog;
use verilog.vl_types.all;
entity xor_testbench is
end xor_testbench;
